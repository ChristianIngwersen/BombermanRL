0.028223230680923896,0.028223230680923896,0.028223230680923896
0.7978101971557853,0.7978101971557853,0.7978101971557853
0.7814789915966386,0.7706770208083233,0.7814147007950696
